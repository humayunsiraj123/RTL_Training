//algo pr =0 ,size [0:2**n-1];
//for i=n-1:to 0;
//   r={pr<<1,a_i}  ;
//  d=r-B;
//  if D<0 so qi =0 ;r =pr
    //else q=1 r=d;
// r= pr;

    
//PR partial remainder  
module full_adder(input a,input b,cin

module div_block(
  input R,
  input B,
  input cin,
  input N,
  output logic PR,
  output logic cout,
  output logic D);
  
              
  
